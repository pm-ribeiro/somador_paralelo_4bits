Somador 4 bits - Concepcao de Circuitos Integrados


* Asterisco indica um COMENTARIO


** Modelo dos transistores
.include ami_035u.mod


** Fonte de alimentação VDD
** Vnome nó+ nó- valor
VDD 1 0 3.3V
VGND GND 0 0V



** Fonte de entrada
** Vnome nó+ nó- PULSE(V1 V2 TD TR TF PW PER)
Vin A1 0 PULSE(0 3.3 0 0.1nS 0.1ns 10ns 20.2ns)
Vin2 A2 0 PULSE(0 3.3 0 0.1nS 0.1ns 20.1ns 40.4ns)
Vin3 A3 0 PULSE(0 3.3 0 0.1nS 0.1ns 40.3ns 80.8ns)
Vin4 A4 0 PULSE(0 3.3 0 0.1nS 0.1ns 80.7ns 170.6ns)
**Vin5 B1 0 PULSE(0 3.3 0 0.1nS 0.1ns 16.8ns 35.2ns)
**Vin6 B2 0 PULSE(0 3.3 0 0.1nS 0.1ns 33.6ns 70.4ns)
**Vin7 B3 0 PULSE(0 3.3 0 0.1nS 0.1ns 67.2ns 140.8ns)
**Vin8 B4 0 PULSE(0 3.3 0 0.1nS 0.1ns 134.4ns 281.6ns)
** Formato de chamada de um transistor MOSFET
** Mnome nó_dreno nó_gate nó_fonte nó_bulk tipo W= L=
.subckt and2 IN IN2 S1 1 GND
M1 OUT IN 1 1 CMOSP W=500u L=0.3u
M2 OUT IN2 1 1 CMOSP W=500u L=0.3u

M3 OUT IN Y 0 CMOSN W=250u L=0.3u
M4 Y IN2 0 0 CMOSN W=250u L=0.3u

X7 OUT S1 1 0 INV
.ends

.subckt or3 A B C S1 1 GND
M1 ADBF A 1 1 CMOSP W=500u L=0.3u
M2 BDCF B ADBF 1 CMOSP W=500u L=0.3u
M3 OUT C BDCF 1 CMOSP W=500u L=0.3u

M4 0 A OUT 0 CMOSN W=250u L=0.3u
M5 0 B OUT 0 CMOSN W=250u L=0.3u
M6 0 C OUT 0 CMOSN W=250u L=0.3u

X7 OUT S1 1 0 INV
.ends

.SUBCKT XOR2 A B SF 1 GND
**inverte a
X1 A AN 1 0 INV
**inverte b
X2 B BN 1 0 INV
**and a e b
X3 AN B S1 1 0 and2
X4 A BN S2 1 0 and2

**or final
M11 ADBF S1 1 1 CMOSP W=500u L=0.3u
M12 OUT S2 ADBF 1 CMOSP W=500u L=0.3u

M14 0 S1 OUT 0 CMOSN W=250u L=0.3u
M15 0 S2 OUT 0 CMOSN W=250u L=0.3u

**inversor
X5 OUT SF 1 0 INV
.ENDS

.SUBCKT INV A SF 1 GND
M17 SF A 1 1 CMOSP W=500u L=0.3u
M18 0 A SF 0 CMOSN W=250u L=0.3u
.ENDS

.subckt SomadorCompleto A B C CARRY SOMA 1 GND
**XOR3
X1 A B SM 1 0 XOR2
X2 SM C SOMA 1 0 XOR2
**Carry
X3 A B S1 1 0 and2
X4 A C S2 1 0 and2
X5 B C S3 1 0 and2
X6 S1 S2 S3 CARRY 1 0 or3
.ENDS

.subckt MS A B CARRY SOMA 1 GND
X1 A B SOMA 1 0 XOR2
X2 A B CARRY 1 0 and2
.ENDS

.subckt Somador4bits A1 A2 A3 A4 B1 B2 B3 B4 S_MS S_SC1 S_SC2 S_SC3 OVER 1 GND
X1 A1 B1 C_MS S_MS 1 0 MS
X2 A2 B2 C_MS C_SC1 S_SC1 1 0 SomadorCompleto
X3 A3 B3 C_SC1 C_SC2 S_SC2 1 0 SomadorCompleto
X4 A4 B4 C_SC2 C_SC3 S_SC3 1 0 SomadorCompleto
X5 C_SC3 C_SC2 OVER 1 0 XOR2
.ENDS
X1 A1 A2 A3 A4 1 1 1 0 S_MS S_SC1 S_SC2 S_SC3 OVER 1 0 Somador4bits

* CAPACITOR DE SAIDA
** Cnome  nó+ nó- valor
C1 S_MS 0 0.10pF
C2 S_SC1 0 0.10pF
C3 S_SC2 0 0.10pF
C4 S_SC3 0 0.10pF
C5 OVER 0 0.1pF


** Analise do transiente
** .tran passo tempo_total
.tran 0.001ns 190ns


** Mostra o grafico
.probe


** Fim da descricao
.end


